// Interface of ham
interface ham_if ();
  logic [7:0] a, b;
  logic [3:0] distance;
endinterface