interface arb_if(input logic clk, rst);
    logic [1:0] r;
    logic [1:0] g;
endinterface //arb_iflogic