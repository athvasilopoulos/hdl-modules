interface bcd_if(input logic clk, rst);
	logic [3:0] ones, tens, hundreds;
endinterface